library verilog;
use verilog.vl_types.all;
entity decoder4to16_vlg_vec_tst is
end decoder4to16_vlg_vec_tst;
