library verilog;
use verilog.vl_types.all;
entity latch2_vlg_vec_tst is
end latch2_vlg_vec_tst;
