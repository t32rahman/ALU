library verilog;
use verilog.vl_types.all;
entity stateMachine_vlg_vec_tst is
end stateMachine_vlg_vec_tst;
